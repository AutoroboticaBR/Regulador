*                                               Revised: Thursday, December 21, 2000
* C:\MEUS DOCUMENTOS\MEUS DOCUMENTOS\REGULADOR.DRevision: 
* 
* 
* 
* 
* 
U1 N00022 N00040 N00025 LM317
R1 N00025 N00040 220R
R2 N00040 N00072 N00072 10K
R3 N00062 N00072 1,5K
J1 N00072 N00019 24v
J2 N00025 N00072 SAIDA
D1 N00019 N00022 1N4007
D2 N00025 N00062 LED
.END
